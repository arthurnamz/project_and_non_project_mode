
`timescale 1ns/1ps


module cpu
#( 
  parameter DATA_WIDTH  = 10,
  parameter MEM_DEPTH  = 8,
  parameter ADDR_WIDTH  = 3
)
( 
   input clk,
   input rstn,
   input start,
   output reg done

);

parameter IDLE = 0;
parameter FETCH = 1;
parameter DEC = 2;
parameter LOAD_OP = 3;
parameter EXEC = 4;
parameter WRITE_BACK = 5;


reg [2:0] state;

// Memory arrays
reg [DATA_WIDTH-1:0] instruction_mem[0:MEM_DEPTH-1];
reg [7:0] data_mem[0:MEM_DEPTH-1];

// Decoded addresses
reg opCode;
reg [2:0] op1;
reg [2:0] op2;
reg [2:0] res;

// Data registers (hold actual values from memory)
reg [7:0] operand1;
reg [7:0] operand2;
reg [7:0] result;

reg [2:0] pc;

// Control signals (generated by combinational block, used by sequential block)
reg pc_inc;
reg pc_reset;

//==================================================================
// SEQUENTIAL LOGIC: State transitions and register/memory updates
//==================================================================
always@(posedge clk) begin
	if(~rstn) begin
		state <= IDLE;
		pc <= 3'd0;
		done <= 1'b0;
		opCode <= 1'b0;
		op1 <= 3'd0;
		op2 <= 3'd0;
		res <= 3'd0;
		operand1 <= 8'd0;
		operand2 <= 8'd0;
		result <= 8'd0;
	end else begin
        // State transitions
        case (state)
            IDLE:   
                if(start)
                    state <= FETCH; 
            FETCH:
                state <= DEC; 
            DEC:
                state <= LOAD_OP;
            LOAD_OP:
                state <= EXEC;
            EXEC:
                state <= WRITE_BACK;
            WRITE_BACK: begin
                if(pc == 3'd7)
                    state <= IDLE;
                else
                    state <= FETCH;
            end
        endcase
        
        // PC update based on control signals
        if(pc_reset)
            pc <= 3'd0;
        else if(pc_inc)
            pc <= pc + 1'b1;
        
        // State-specific operations
        case(state)
            DEC: begin
                opCode <= instruction_mem[pc][0];
                op1 <= instruction_mem[pc][3:1];
                op2 <= instruction_mem[pc][6:4];
                res <= instruction_mem[pc][9:7];
            end
            
            LOAD_OP: begin
                operand1 <= data_mem[op1];
                operand2 <= data_mem[op2];
            end
            
            EXEC: begin
                if(opCode == 1'b0)
                    result <= operand1 + operand2;
                else
                    result <= ~operand1;
            end
            
            WRITE_BACK: begin
                data_mem[res] <= result;
                if(pc == 3'd7)
                    done <= 1'b1;
                else
                    done <= 1'b0;
            end
        endcase
    end
end	

//==================================================================
// COMBINATIONAL LOGIC: Generate control signals based on state
//==================================================================
always @(*) begin
    // Default values
    pc_inc = 1'b0;
    pc_reset = 1'b0;
    
	case(state)
        IDLE: begin
            pc_reset = 1'b1;
        end
        
        WRITE_BACK: begin
            pc_inc = 1'b1;
        end
	endcase
end


endmodule
